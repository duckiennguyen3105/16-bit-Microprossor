LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY mux3_1 IS
PORT ( X,Y : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Z : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		S : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		M : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END  mux3_1;

ARCHITECTURE Behavior OF mux3_1 IS
BEGIN
	PROCESS(S,X,Y,Z)
	BEGIN
		CASE S IS
			WHEN "00" => M <= Y;
			WHEN "01" => M <="00000000" & Z;
			WHEN "10" => M <= X;
			WHEN OTHERS => NULL;
		END CASE;
	END PROCESS;

END Behavior;

